`ifndef __INSTRUCTIONDECODE__
`define __INSTRUCTIONDECODE__

module instructionDecode
(
  input [31:0] instruction,

  //outputs for each possible instruction 
  //outputs for rd, rs1, rs2, and immediates
  //outputs for if rd, rs1, rs2, and immediates are used/valid
);

`endif
